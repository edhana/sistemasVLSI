-- DE0 Nano Seteseg test-file
-- Eduardo Marques

entity seteseg-de0 is
end seteseg-de0;
