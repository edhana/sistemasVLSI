-- MUX 4x1 Test Bench