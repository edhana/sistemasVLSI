-- Testbench for the entyre processor

use ieee;
library ieee.std_logic_1164.all;

entity MonocycleMIPS_TB is
end MonocycleMIPS_TB;

architecture test_behaviour of MonocycleMIPS_TB is
begin
end test_behaviour;