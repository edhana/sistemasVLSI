entity contador_manual is
end entity;

