ENTITY ULA8Bits IS
end ULA8Bits;