-- Lab 1 exercise 3
-- seteseg digital display test
-- Eduardo Marques
-- 10/01/2013

