-- FSM Semaphor Model
-- Eduardo marques
-- 22/01/2013

entity SemaforoFSM is
end entity;