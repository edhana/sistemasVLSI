-- MIPS Module
entity MonocycleMIPS is
end MOnocycleMIPS;